module inverse(y, x);
	input [4:0] x;
	output [4:0] y;
	reg [4:0] y;
	always @ (x)
	case (x) 
		1: y = 1; 
		2: y = 18; 
		4: y = 9; 
		8: y = 22; 
		16: y = 11; 
		5: y = 23; 
		10: y = 25; 
		20: y = 30; 
		13: y = 15; 
		26: y = 21; 
		17: y = 24; 
		7: y = 12; 
		14: y = 6; 
		28: y = 3; 
		29: y = 19; 
		31: y = 27; 
		27: y = 31; 
		19: y = 29; 
		3: y = 28; 
		6: y = 14; 
		12: y = 7; 
		24: y = 17; 
		21: y = 26; 
		15: y = 13; 
		30: y = 20; 
		25: y = 10; 
		23: y = 5; 
		11: y = 16; 
		22: y = 8; 
		9: y = 4; 
		18: y = 2; 
	endcase
endmodule