module BUFFER (OUT,IN);
    input IN;
    output OUT;
        buf (OUT, IN);
endmodule