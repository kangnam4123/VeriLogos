module vd30ca9_vb2eccd (
 output q
);
 assign q = 1'b0;
endmodule