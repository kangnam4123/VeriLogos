module mbuf (
	   input a,
	   output q
	   );
   assign 	  q = a;
endmodule