module vcdce79_v9a2a06 (
 input i1,
 input [3:0] i0,
 output [4:0] o
);
 assign o = {i1, i0};
endmodule