module AND2_3 (
	input A, B,
	output Y
);
	assign Y = A & B;
endmodule