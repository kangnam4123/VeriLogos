module MuxN_14(
  input  [31:0] io_ins_0,
  output [31:0] io_out
);
  wire [31:0] _GEN_0;
  assign io_out = _GEN_0;
  assign _GEN_0 = io_ins_0;
endmodule