module TIEHHD (Z);
output Z ;
   buf (Z, 1'B1);
endmodule