module vd12401_vf4938a (
 input a,
 input b,
 output c
);
 assign c = a ^ b;
endmodule