module abc9_test024_sub(input [1:0] i, output [1:0] o);
assign o = i;
endmodule