module Arbiter_8(
  output  io_in_0_ready,
  input   io_out_ready
);
  assign io_in_0_ready = io_out_ready; 
endmodule