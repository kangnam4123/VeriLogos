module abc9_test003(input [1:0] a, output [1:0] o);
assign o = a;
endmodule