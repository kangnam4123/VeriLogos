module twentynm_io_ibuf (output o, input i, input ibar);
   assign ibar = ibar;
   assign o    = i;
endmodule