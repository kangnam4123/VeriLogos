module NV_BLKBOX_SRC0 (
  Y
 );
output Y ;
assign Y = 1'b0;
endmodule