module BUFF_2 (o, i);
    output o;
    input i;
    assign o = i;
endmodule