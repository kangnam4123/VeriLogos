module JAND2B(A1, A2, O);
input   A1;
input   A2;
output  O;
and g0(O, A1, A2);
endmodule