module v4c802f_v465065 #(
 parameter VALUE = 0
) (
 output [23:0] k
);
 assign k = VALUE;
endmodule