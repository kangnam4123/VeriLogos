module SyncReset0 (
		   IN_RST_N,
		   OUT_RST_N
		   );
   input   IN_RST_N ;
   output  OUT_RST_N ;
   assign  OUT_RST_N = IN_RST_N ;
endmodule