module JCINVA1(A, O);
input   A;
output  O;
not g0(O, A);
endmodule