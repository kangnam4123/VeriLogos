module test_19(p);
   output p;
   assign q = 1; 
   assign p = q;
endmodule