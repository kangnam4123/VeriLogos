module f6 (a, b, clk, q);
   input  [2:0] a;
   input [2:0] 	b;
   input 	clk;
   output 	q;
   reg 		out;
   function func6;
      reg 	result;
      input [5:0] src;
      begin
	 if (src[5:0] == 6'b011011) begin
	    result = 1'b1;
	 end
	 else begin
	    result = 1'b0;
	 end
	 func6 = result;
      end
   endfunction
   wire [5:0] w6 = {a, b};
   always @(posedge clk) begin
      out <= func6(w6);
   end
   assign q = out;
endmodule