module hardcaml_lib_gnd
(
    output o
);
    assign o = 1'b0;
endmodule