module f1_TECH_AND18(input [17:0] in, output out);
assign out = &in;
endmodule