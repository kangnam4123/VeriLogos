module feedx1 (Z, A);
  output Z;
  input A;
  assign Z = A;
endmodule