module logic_1(output a);
    assign a = 1;
endmodule