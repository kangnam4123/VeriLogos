module r_USBPD_REV_VER_LOW(output wire [7:0] reg_0x08);
	assign reg_0x08=8'h00;
endmodule