module cp_u4l(output wire logic unsigned [11:0] dst,
              input  wire logic unsigned [11:0] src);
  assign dst = src;
endmodule