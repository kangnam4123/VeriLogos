module my_and_1 (out,a,b);
input a,b;
output out;
and u0 (out,a,b);
endmodule