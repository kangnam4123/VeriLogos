module a (input i, output oa);
   assign i = 1'b1;
   assign oa = i;
endmodule