module One;
   wire one = 1'b1;
endmodule