module MJNOR8C(A1, A2, A3, A4, A5, A6, A7, A8, O);
input   A1;
input   A2;
input   A3;
input   A4;
input   A5;
input   A6;
input   A7;
input   A8;
output  O;
nor g0(O, A1, A2, A3, A4, A5, A6, A7, A8);
endmodule