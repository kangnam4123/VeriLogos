module lab5iram1B(CLK, RESET, ADDR, Q);
  input         CLK;
  input         RESET;
  input  [7:0]  ADDR;
  output [15:0] Q;
  reg    [15:0] mem[0:127]; 
  wire   [6:0]  saddr;
  integer       i;
  assign saddr = ADDR[7:1];
  assign Q = mem[saddr];
  always @(posedge CLK) begin
    if(RESET) begin
      mem[0]  <= 16'b1111000000000001; 
      mem[1]  <= 16'b0101000101111111; 
      mem[2]  <= 16'b0010101001111010; 
      mem[3]  <= 16'b0010101010111011; 
      mem[4]  <= 16'b0100101001000000; 
      mem[5]  <= 16'b0100101010111111; 
      mem[6]  <= 16'b0110010011000001; 
      mem[7]  <= 16'b1111000011011001; 
      mem[8]  <= 16'b1111001011011101; 
      mem[9]  <= 16'b1111000011100000; 
      mem[10]  <= 16'b1111001000001100; 
      mem[11]  <= 16'b1111010000010011; 
      mem[12]  <= 16'b0110010011000001; 
      mem[13]  <= 16'b1111000011011001; 
      mem[14]  <= 16'b1111001011011101; 
      mem[15]  <= 16'b1111100011100000; 
      mem[16]  <= 16'b1111001000001100; 
      mem[17]  <= 16'b1111010000010011; 
      mem[18]  <= 16'b0110010011000001; 
      mem[19]  <= 16'b1111000011011001; 
      mem[20]  <= 16'b1111001011011101; 
      mem[21]  <= 16'b1111100011100000; 
      mem[22]  <= 16'b1111001000001100; 
      mem[23]  <= 16'b1111010000010011; 
      mem[24]  <= 16'b0110010011000001; 
      mem[25]  <= 16'b1111000011011001; 
      mem[26]  <= 16'b1111001011011101; 
      mem[27]  <= 16'b1111100011100000; 
      mem[28]  <= 16'b0100101100111110; 
      mem[29]  <= 16'b0010101100111100; 
      mem[30]  <= 16'b0100101100111101; 
      for(i = 31; i < 128; i = i + 1) begin
        mem[i] <= 16'b0000000000000000;
      end
    end
  end
endmodule