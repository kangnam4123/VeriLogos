module inv_3(o,i);
input i;
output o;
assign o = ~i;
endmodule