module GP_VDD(output OUT);
       assign OUT = 1;
endmodule