module GSR_3(output GSR);
    assign GSR = 1'b1;
endmodule