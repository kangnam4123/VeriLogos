module r_DEVICE_ID_LOW(output wire [7:0] reg_0x04);
	assign reg_0x04=8'h00;
endmodule