module r_PD_INTERFACE_REV_LOW(output wire [7:0] reg_0x0A);
	assign reg_0x0A=8'h00;
endmodule