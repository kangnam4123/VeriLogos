module sysgen_constant_737c6ebc01 (
  output [(4 - 1):0] op,
  input clk,
  input ce,
  input clr);
  assign op = 4'b1111;
endmodule