module alpha_3 (
   toggle_up,
   clk, toggle, cyc_copy
   );
   input clk;
   input toggle;
   input [7:0] cyc_copy;
   reg 	       toggle_internal;
   output reg  toggle_up;
   always @ (posedge clk) begin
      toggle_internal <= toggle;
      toggle_up       <= toggle;
   end
endmodule