module MJNOR2B1(A1, A2, O);
input   A1;
input   A2;
output  O;
nor g0(O, A1, A2);
endmodule