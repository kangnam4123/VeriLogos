module bug34649 (name);
       output reg name = 0;
endmodule