module bug27039;
   integer i;
endmodule