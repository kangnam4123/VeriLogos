module nios_solo_nios2_gen2_0_cpu_nios2_oci_pib (
                                                   tr_data
                                                )
;
  output  [ 35: 0] tr_data;
  wire    [ 35: 0] tr_data;
  assign tr_data = 0;
endmodule