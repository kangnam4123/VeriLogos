module CONNECTNET(IN, OUT);
output OUT;
input IN;
assign OUT = IN;
endmodule