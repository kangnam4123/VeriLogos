module v651fa3_v465065 #(
 parameter VALUE = 0
) (
 output [15:0] k
);
 assign k = VALUE;
endmodule