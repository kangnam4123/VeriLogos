module lcd (clk, lcd_rs, lcd_rw, lcd_e, lcd_0, lcd_1, lcd_2, lcd_3, lcd_4, lcd_5, lcd_6, lcd_7);
                    parameter       k = 18;
   input           clk;        
                    reg   [k+8-1:0] count=0;
                    reg             lcd_busy=1;
                    reg             lcd_stb;
                    reg       [5:0] lcd_code;
                    reg       [6:0] lcd_stuff;
   output reg      lcd_rs;
   output reg      lcd_rw;
   output reg      lcd_7;
   output reg      lcd_6;
   output reg      lcd_5;
   output reg      lcd_4; 
     output reg      lcd_3;
     output reg      lcd_2;
     output reg      lcd_1;
     output reg      lcd_0;
   output reg      lcd_e;
  always @ (posedge clk) begin
    count  <= count + 1;
 lcd_0 <= 0;
 lcd_1 <= 0;
 lcd_2 <= 0;
 lcd_3 <= 0;
    case (count[k+7:k+2])
       0: lcd_code <= 6'h03;        
       1: lcd_code <= 6'h03;
       2: lcd_code <= 6'h03;
       3: lcd_code <= 6'h02;
       4: lcd_code <= 6'h02;        
       5: lcd_code <= 6'h08;
       6: lcd_code <= 6'h00;        
       7: lcd_code <= 6'h06;
       8: lcd_code <= 6'h00;        
       9: lcd_code <= 6'h0C;
      10: lcd_code <= 6'h00;        
      11: lcd_code <= 6'h01;
		12: lcd_code <= 6'h22;        
      13: lcd_code <= 6'h2A;
      14: lcd_code <= 6'h22;        
      15: lcd_code <= 6'h20;
      16: lcd_code <= 6'h24;        
      17: lcd_code <= 6'h23;
      18: lcd_code <= 6'h24;        
      19: lcd_code <= 6'h2F;
      20: lcd_code <= 6'h24;        
      21: lcd_code <= 6'h2C;
      22: lcd_code <= 6'h24;        
      23: lcd_code <= 6'h25;
      24: lcd_code <= 6'h24;        
      25: lcd_code <= 6'h23;
      26: lcd_code <= 6'h24;        
      27: lcd_code <= 6'h2F;
      28: lcd_code <= 6'h25;        
      29: lcd_code <= 6'h26;
      30: lcd_code <= 6'h24;        
      31: lcd_code <= 6'h29;
      32: lcd_code <= 6'h25;        
      33: lcd_code <= 6'h23;
      34: lcd_code <= 6'h24;        
      35: lcd_code <= 6'h29;
		36: lcd_code <= 6'h24;        
      37: lcd_code <= 6'h2F;
		38: lcd_code <= 6'h24;        
      39: lcd_code <= 6'h2E;
		40: lcd_code <= 6'h22;        
      41: lcd_code <= 6'h20;
		42: lcd_code <= 6'h22;        
      43: lcd_code <= 6'h2A;
      default: lcd_code <= 6'h10;
    endcase
  if (lcd_rw)                     
    lcd_busy <= 0;                
    lcd_stb <= ^count[k+1:k+0] & ~lcd_rw & lcd_busy;  
    lcd_stuff <= {lcd_stb,lcd_code};
    {lcd_e,lcd_rs,lcd_rw,lcd_7,lcd_6,lcd_5,lcd_4} <= lcd_stuff;
  end
endmodule