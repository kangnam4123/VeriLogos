module NV_BLKBOX_BUFFER (
  Y
 ,A
 );
output Y ;
input A ;
assign Y = A;
endmodule