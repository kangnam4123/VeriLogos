module InstruMemory 
#(parameter DATA_WIDTH = 32, parameter ADDR_WIDTH = 32)
(
	input [(DATA_WIDTH-1):0] data,
	input [(ADDR_WIDTH-1):0] addr,
	input [3:0] we, 
	input clk,
	output [(DATA_WIDTH-1):0] q
);
	reg [DATA_WIDTH-1:0] ram[2**(ADDR_WIDTH - 22) - 1:0];
	reg [ADDR_WIDTH-1:0] addr_reg;
initial
begin
ram[0] = 32'b000000_01001_01010_00011_00000_100000;
ram[1] = 32'b000000_01001_01100_00100_00000_100010;
ram[2] = 32'b000000_11111_00100_00101_00000_100010;
ram[3] = 32'b000000_00101_00001_00011_00000_100000;
ram[4] = 32'b000000_00100_00001_00101_00000_100011;
ram[5] = 32'b000000_00010_00101_00101_00000_000111;
ram[6] = 32'b000000_00010_01001_00101_00010_000010;
ram[7] = 32'b000000_01010_01001_00101_00000_101011;
ram[8] = {16'b001000_00101_00101,16'h789a};
ram[9] = {16'b001000_11111_00101,16'h7abc};
ram[10] = {16'b001001_11111_00101,16'h7abc};
ram[11] = {16'b001001_00101_00101,16'h789a};
ram[12] = {16'b001111_00000_00101,16'h789a};
ram[13] = {16'b001110_11111_00101,16'habcd};
ram[14] = 32'b011100_01011_00010_00101_00000_100001;
ram[15] = 32'b011100_01010_00010_00101_00000_100000;
ram[16] = {16'b001010_00101_00101,16'habcd};
ram[17] = 32'b011111_00000_01101_00110_10000_100000;
ram[18] = {16'b101011_00000_01001,16'd512};
ram[19] = {16'b101010_00000_11111,16'd256};
ram[20] = {16'b100011_00000_00011,16'd512};
ram[21] = {16'b100010_00000_00011,16'd513};
ram[22] = {16'b100010_00000_00011,16'd514};
ram[23] = {16'b100010_00000_00011,16'd515};
ram[24] = {16'b100110_00000_00011,16'd513};
ram[25] = {16'b100110_00000_00011,16'd514};
ram[26] = {16'b100110_00000_00011,16'd515};
ram[27] = 32'b000000_01001_00011_00011_00000_100000;
ram[28] = {16'b101010_00000_11111,16'd513};
ram[29] = {16'b101010_00000_11111,16'd514};
ram[30] = {16'b101010_00000_11111,16'd515};
ram[31] = {16'b101110_00000_11111,16'd513};
ram[32] = {16'b101110_00000_11111,16'd514};
ram[33] = {16'b101110_00000_11111,16'd515};
ram[34] = {16'b000001_00001_10001,16'h0006};
ram[35] = {6'b000010,2'b0,24'h0};
ram[41] = {16'b000001_11110_00001,16'h0001};
ram[42] = {6'b000010,2'b0,24'h0};
end
	always @ (negedge clk)
	begin
		if (we[0] == 1'b1)
			ram[addr[9:2]][7:0] <= data[7:0];
		if (we[1] == 1'b1)
			ram[addr[9:2]][15:8] <= data[15:8];
		if (we[2] == 1'b1)
			ram[addr[9:2]][23:16] <= data[23:16];
		if (we[3] == 1'b1)
			ram[addr[9:2]][31:24] <= data[31:24];
	end
	assign q = ram[addr[9:2]];
endmodule