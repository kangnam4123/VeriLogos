module v9b9118_v465065 #(
 parameter VALUE = 0
) (
 output [3:0] k
);
 assign k = VALUE;
endmodule