module SUB1(input in1, in2, cin, output out, cout);
assign {cout, out} = in1 - in2 - cin;
endmodule