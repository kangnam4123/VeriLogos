module N1Z001( O );     
    output  O;
assign O = 1'b1;
endmodule