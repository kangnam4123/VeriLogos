module SYN_IBUF_1(input I, output O);
  assign O = I;
endmodule