module f3_test_1(in, out);
input wire in;
output  out;
assign out = (in+in);
assign out = 74;
endmodule