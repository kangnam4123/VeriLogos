module f12_test(input in, output out);
assign out = in;
endmodule