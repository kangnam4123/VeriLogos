module sysgen_constant_bd840882a6 (
  output [(32 - 1):0] op,
  input clk,
  input ce,
  input clr);
  assign op = 32'b00000100100000000000000000000000;
endmodule