module ident(
	     input  i_ident,
	     output o_ident
	     );
   assign o_ident = i_ident;
endmodule