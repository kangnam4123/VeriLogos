module sub_25;
   integer inside_sub_a = 1;
endmodule