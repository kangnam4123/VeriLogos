module BUFF (
	input A,
	output Y
);
	assign Y = A;
endmodule