module sky130_fd_sc_hvl__lsbufhv2hv_hl_1 (
    X,
    A
);
    output X;
    input  A;
    buf buf0 (X     , A              );
endmodule