module SYN_OBUF_1(input I, output O);
  assign O = I;
endmodule