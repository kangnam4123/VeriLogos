module BUFG_6(I, O);
    input I;
    output O;
    assign O = I;
endmodule