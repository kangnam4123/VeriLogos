module Gi(input A, input B, output G);
	assign G = A&B;
endmodule