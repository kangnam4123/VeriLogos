module buff_1 (
    output Q,
    input  A
);
  assign Q = A;
endmodule