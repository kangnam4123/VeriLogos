module r_DEVICE_ID_HIGH(output wire [7:0] reg_0x05);
	assign reg_0x05=8'h00;
endmodule