module f1_test_5(input in, output out);
assign out = in;
endmodule