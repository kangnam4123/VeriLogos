module m_2 (x);
   output x;
   reg	  x;
endmodule