module BUF_1(DATA, RESULT);
input DATA;
output RESULT;
assign RESULT = DATA;
endmodule