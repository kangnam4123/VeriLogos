module BUFG_2(I,O);
input I;
output O;
assign #1 O=I;
endmodule