module INVX4(A, Y);
input A;
output Y;
not(Y, A);
endmodule