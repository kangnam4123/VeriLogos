module mgc_io_sync (ld, lz);
    input  ld;
    output lz;
    assign lz = ld;
endmodule