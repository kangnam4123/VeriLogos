module add_sub27(add, opa, opb, sum, co);
input		add;
input	[26:0]	opa, opb;
output	[26:0]	sum;
output		co;
assign {co, sum} = add ? (opa + opb) : (opa - opb);
endmodule