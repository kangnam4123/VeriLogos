module CPE_base (x,y,Int_pel,out);
	input [3:0] x;	
	input [3:0] y;	
	input [7:0] Int_pel;
	output [13:0] out;
	wire [10:0] sum_x3;
	wire [9:0] sum_x2;
	wire [8:0] sum_x1;
	wire [7:0] sum_x0;
	wire [10:0] sum_x;
	wire [13:0] sum_y3;
	wire [12:0] sum_y2;
	wire [11:0] sum_y1;
	wire [10:0] sum_y0;
	assign sum_x3 = (x[3] == 1'b1)? {Int_pel,3'b0}:0;
	assign sum_x2 = (x[2] == 1'b1)? {Int_pel,2'b0}:0;
	assign sum_x1 = (x[1] == 1'b1)? {Int_pel,1'b0}:0;
	assign sum_x0 = (x[0] == 1'b1)? Int_pel:0; 
	assign sum_x = (sum_x3 + sum_x2) + (sum_x1 + sum_x0);
	assign sum_y3 = (y[3] == 1'b1)? {sum_x,3'b0}:0;
	assign sum_y2 = (y[2] == 1'b1)? {sum_x,2'b0}:0;
	assign sum_y1 = (y[1] == 1'b1)? {sum_x,1'b0}:0;
	assign sum_y0 = (y[0] == 1'b1)? sum_x:0; 
	assign out = (sum_y3 + sum_y2) + (sum_y1 + sum_y0);
endmodule