module MSCINVD3 (O,A);
    output O;
    input A;
        not             U_1     ( O , A);
endmodule