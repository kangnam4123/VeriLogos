module ma_1(x);
  output [3:0] x;
  parameter P = 4'd5;
  assign x = P;
endmodule