module r_PRODUCT_ID_HIGH(output wire [7:0] reg_0x03);
	assign reg_0x03=8'h00;
endmodule