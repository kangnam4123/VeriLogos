module LUT_SHIFT_1 #(parameter P = 32, parameter D = 5) ( 
input wire CLK, 
input wire EN_ROM1,
input wire [D-1:0] ADRS,
output reg [P-1:0] O_D
);
always @(posedge CLK)
      if (EN_ROM1)
         case (ADRS)
            5'b00000: O_D <= 32'b00111111011111110000000000000000;
            5'b00001: O_D <= 32'b00111111011111100000000000000000;
            5'b00010: O_D <= 32'b00111111011111000000000000000000;
            5'b00011: O_D <= 32'b00111111011110000000000000000000;
            5'b00100: O_D <= 32'b00111111011100000000000000000000;
            5'b00101: O_D <= 32'b00111111011000000000000000000000;
            5'b00110: O_D <= 32'b00111111010000000000000000000000;
            5'b00111: O_D <= 32'b00111111000000000000000000000000;
            5'b01000: O_D <= 32'b00111110100000000000000000000000;
            5'b01001: O_D <= 32'b00111110000000000000000000000000;
            5'b01010: O_D <= 32'b00111101100000000000000000000000;
            5'b01011: O_D <= 32'b00111101100000000000000000000000;
            5'b01100: O_D <= 32'b00111101000000000000000000000000;
            5'b01101: O_D <= 32'b00111100100000000000000000000000;
            5'b01110: O_D <= 32'b00111100000000000000000000000000;
            5'b01111: O_D <= 32'b00111100000000000000000000000000;
            5'b10000: O_D <= 32'b00111011100000000000000000000000;
            5'b10001: O_D <= 32'b00111011000000000000000000000000;
            5'b10010: O_D <= 32'b00111010100000000000000000000000;
            5'b10011: O_D <= 32'b00111010000000000000000000000000;
            5'b10100: O_D <= 32'b00111010000000000000000000000000;
            5'b10101: O_D <= 32'b00111001100000000000000000000000;
            5'b10110: O_D <= 32'b00111001000000000000000000000000;
            5'b10111: O_D <= 32'b00111000011111111111111111111110;
            5'b11000: O_D <= 32'b00111000011111111111111111111110;
            5'b11001: O_D <= 32'b00110111111111111111111111111100;
            5'b11010: O_D <= 32'b00110111011111111111111111110110;
            5'b11011: O_D <= 32'b00110111011111111111111111110110;
            5'b11100: O_D <= 32'b00110110111111111111111111110110;
            5'b11101: O_D <= 32'b00110110011111111111111111100000;
            5'b11110: O_D <= 32'b00110110011111111111111111100000;
            5'b11111: O_D <= 32'b00110101111111111111111110110100;
            default:  O_D <= 32'b00000000000000000000000000000000;
        endcase
endmodule