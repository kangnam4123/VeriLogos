module altera_up_avalon_video_dma_ctrl_addr_trans (
	clk,
	reset,
	slave_address,
	slave_byteenable,
	slave_read,
	slave_write,
	slave_writedata,
	master_readdata,
	master_waitrequest,
	slave_readdata,
	slave_waitrequest,
	master_address,
	master_byteenable,
	master_read,
	master_write,
	master_writedata
);
parameter ADDRESS_TRANSLATION_MASK	= 32'hC0000000;
input					clk;
input					reset;
input			[ 1: 0]	slave_address;
input			[ 3: 0]	slave_byteenable;
input					slave_read;
input					slave_write;
input			[31: 0]	slave_writedata;
input			[31: 0]	master_readdata;
input					master_waitrequest;
output			[31: 0]	slave_readdata;
output					slave_waitrequest;
output			[ 1: 0]	master_address;
output			[ 3: 0]	master_byteenable;
output					master_read;
output					master_write;
output			[31: 0]	master_writedata;
assign slave_readdata		= (slave_address[1] == 1'b0) ? 
								master_readdata | ADDRESS_TRANSLATION_MASK :
								master_readdata;
assign slave_waitrequest	= master_waitrequest;
assign master_address		= slave_address;
assign master_byteenable	= slave_byteenable;
assign master_read			= slave_read;
assign master_write			= slave_write;
assign master_writedata		= (slave_address[1] == 1'b0) ?
								slave_writedata & ~ADDRESS_TRANSLATION_MASK :
								slave_writedata;
endmodule