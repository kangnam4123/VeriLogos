module xor3(input a ,input b,input c,output x);
   assign x=a^b^c;
endmodule