module IV2(A,  Z);
  input A;
  output Z;
  assign Z = ~A;
endmodule