module clb_l (input clk, input [15:0] din, output [15:0] dout);
	assign dout = 0;
endmodule