module hardcaml_lib_z
(
    output o
);
    assign o = 1'bz;
endmodule