module INV_8(input A, output Z);
	assign Z = !A;
endmodule