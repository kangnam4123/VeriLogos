module bw_io_dtl_rcv_dc (
  so, 
  pad, ref, vddo
  );
  output	so;
  input		pad;
  input		ref;
  input		vddo;
  assign so = pad ;
  endmodule