module sysgen_constant_9243789fee (
  output [(9 - 1):0] op,
  input clk,
  input ce,
  input clr);
  assign op = 9'b111111111;
endmodule