module v6b14d5_v465065 #(
 parameter VALUE = 0
) (
 output k
);
 assign k = VALUE;
endmodule