module r_FAULT_CONTROL(output reg [7:0] reg_0x1B, input wire reset, input wire wenb, input wire [7:0] in_data, input wire clk);
	always@(posedge clk)
	begin
		if(reset==0) begin
			if(wenb==0)
				reg_0x1B<=in_data;
			else
				reg_0x1B<=reg_0x1B;
		end
		else
			reg_0x1B<=8'h00;
	end
endmodule