module zero(
	output zero);
 	
	assign zero = 1'b0;
	
endmodule