module abc9_test007_sub(input a, output b);
assign b = a;
endmodule