module NV_BLKBOX_SRC0_X(
Y
);
output Y;
assign Y = 1'b0;
endmodule