module thirtytwobitsubtractor(a,b,carryout,s,carryin); 
input [31:0] a,b;
output [31:0] s;
input carryin;
output carryout;
wire [31:0] m;
xor X0(m[0],b[0],1);
xor X1(m[1],b[1],1);
xor X2(m[2],b[2],1);
xor X3(m[3],b[3],1);
xor X4(m[4],b[4],1);
xor X5(m[5],b[5],1);
xor X6(m[6],b[6],1);
xor X7(m[7],b[7],1);
xor X8(m[8],b[8],1);
xor X9(m[9],b[9],1);
xor X10(m[10],b[10],1);
xor X11(m[11],b[11],1);
xor X12(m[12],b[12],1);
xor X13(m[13],b[13],1);
xor X14(m[14],b[14],1);
xor X15(m[15],b[15],1);
xor X16(m[16],b[16],1);
xor X17(m[17],b[17],1);
xor X18(m[18],b[18],1);
xor X19(m[19],b[19],1);
xor X20(m[20],b[20],1);
xor X21(m[21],b[21],1);
xor X22(m[22],b[22],1);
xor X23(m[23],b[23],1);
xor X24(m[24],b[24],1);
xor X25(m[25],b[25],1);
xor X26(m[26],b[26],1);
xor X27(m[27],b[27],1);
xor X28(m[28],b[28],1);
xor X29(m[29],b[29],1);
xor X30(m[30],b[30],1);
xor X31(m[31],b[31],1);
endmodule