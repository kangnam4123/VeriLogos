module GeneratorUnsigned2(out);
	output wire [1:0] out;
	assign out = 2;
endmodule