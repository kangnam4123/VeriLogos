module sysgen_constant_b4741603e8 (
  output [(32 - 1):0] op,
  input clk,
  input ce,
  input clr);
  assign op = 32'b00000111111111110000000000000000;
endmodule