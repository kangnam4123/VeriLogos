module abc9_test002(input [1:0] a, output o);
assign o = a[1];
endmodule