module foo_9(a);
   output a;
   wire a = 1'b1 ;
endmodule