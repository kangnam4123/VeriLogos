module i2c_test02(clk, slave_wait, clk_cnt, cmd, cmd_stop, cnt);
	input clk, slave_wait, clk_cnt;
	input cmd;
	output reg cmd_stop;
	reg clk_en;
	output reg [15:0] cnt;
	always @(posedge clk)
	  if (~|cnt)
	    if (~slave_wait)
	      begin
	          cnt    <= #1 clk_cnt;
	          clk_en <= #1 1'b1;
	      end
	    else
	      begin
	          cnt    <= #1 cnt;
	          clk_en <= #1 1'b0;
	      end
	  else
	    begin
                cnt    <= #1 cnt - 16'h1;
	        clk_en <= #1 1'b0;
	    end
	always @(posedge clk)
	  if (clk_en)
	    cmd_stop <= #1 cmd;
endmodule