module incif_wrapuint8_127_incnil(input CLK, input CE, input [8:0] process_input, output [7:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [7:0] unnamedcast394USEDMULTIPLEcast;assign unnamedcast394USEDMULTIPLEcast = (process_input[7:0]); 
  assign process_output = (((process_input[8]))?((({(unnamedcast394USEDMULTIPLEcast==(8'd127))})?((8'd0)):({(unnamedcast394USEDMULTIPLEcast+(8'd1))}))):(unnamedcast394USEDMULTIPLEcast));
endmodule