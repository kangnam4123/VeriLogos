module bw_io_dtl_vref (
   vref_impctl, vddo
   );
   output        vref_impctl;
   input         vddo;              
assign vref_impctl = 1'b1;
endmodule