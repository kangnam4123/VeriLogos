module ACINVF(A, O);
input   A;
output  O;
not g0(O, A);
endmodule