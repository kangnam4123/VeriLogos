module sub_15;
   reg subsig1 ;
   reg subsig2 ;
endmodule