module mod4 (ident1,out1);
input  [31:0]  ident1;
output [31:0]  out1;
wire [31:0] out1 = ident1;
endmodule