module ChildB(input A, output Y);
  assign Y = A;
endmodule