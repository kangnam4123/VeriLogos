module OR2D1 (
  A1
 ,A2
 ,Z
 );
input A1 ;
input A2 ;
output Z ;
assign Z = A1 | A2;
endmodule