module JBUFNAD(B, A, O);
input   B;
input   A;
output  O;
buf g0(O, B);
endmodule