module dp_mux2es (dout, in0, in1, sel) ;
parameter SIZE = 1;
output 	[SIZE-1:0] 	dout;
input	[SIZE-1:0]	in0;
input	[SIZE-1:0]	in1;
input			sel;
reg	[SIZE-1:0]	dout ;
always @ (sel or in0 or in1)
 begin
	   case (sel)
	     1'b1: dout = in1 ; 
	     1'b0: dout = in0;
	     default: 
         begin
            if (in0 == in1) begin
               dout = in0;
            end
            else
              dout = {SIZE{1'bx}};
         end
	   endcase 
 end
endmodule