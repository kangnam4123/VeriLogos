module cycloneive_io_ibuf_1
  (output o, input i, input ibar);
   assign ibar = ibar;
   assign o    = i;
endmodule