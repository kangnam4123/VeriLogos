module VCC_2 (output V);
   assign V = 1'b1;
endmodule