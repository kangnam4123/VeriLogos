module cp_s4(output wire logic signed [7:0] dst,
             input  wire logic signed [7:0] src);
  assign dst = src;
endmodule