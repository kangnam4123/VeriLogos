module f6_test_3(input in, output out);
assign out = in;
endmodule