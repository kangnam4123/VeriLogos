module NameA ();
parameter ident0 = 12;
parameter ident1 = 20 ;
wire [31:0] value0 = ident0;
wire [31:0] value1 = ident1;
endmodule