module s05;
  integer global; initial global = 1;
endmodule