module XORCY(output O, input CI, LI);
  assign O = CI ^ LI;
endmodule