module OBUF_4(output O, input I);
	assign O = I;
endmodule