module bw_io_ic_filter(
    torcvr,
   topad,
   vddo );
output  torcvr;
input   topad;
input   vddo;
assign torcvr = topad ;
endmodule