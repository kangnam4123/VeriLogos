module NBUFFX8_1 (INP,Z);
	input INP;
	output Z;
assign Z = INP;
endmodule