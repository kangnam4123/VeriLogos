module clock_pkg();
   wire int_clk;
endmodule