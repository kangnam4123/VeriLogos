module incif_wrapuint16_323_incnil(input CLK, input CE, input [16:0] process_input, output [15:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] unnamedcast3810USEDMULTIPLEcast;assign unnamedcast3810USEDMULTIPLEcast = (process_input[15:0]); 
  assign process_output = (((process_input[16]))?((({(unnamedcast3810USEDMULTIPLEcast==(16'd323))})?((16'd0)):({(unnamedcast3810USEDMULTIPLEcast+(16'd1))}))):(unnamedcast3810USEDMULTIPLEcast));
endmodule