module GP_IBUF(input IN, output OUT);
	assign OUT = IN;
endmodule