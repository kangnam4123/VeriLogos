module cn1 (out, in1);
input in1 ;
output out ;
   assign out = in1;
endmodule