module va5ad63_v465065 #(
 parameter VALUE = 0
) (
 output [5:0] k
);
 assign k = VALUE;
endmodule