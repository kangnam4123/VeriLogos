module abc9_test004(input [1:0] a, output o);
assign o = ^a;
endmodule