module BUF_2 (input in, output out);
assign out = in;
endmodule