module one (a);
   input a;
   reg x;
endmodule