module GeneratorSigned2(out);
	output wire signed [1:0] out;
	assign out = 2;
endmodule