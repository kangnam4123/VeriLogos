module sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_3 (
    X,
    A
);
    output X;
    input  A;
    buf buf0 (X     , A              );
endmodule