module INV_14(input in, output out);
assign out = ~in;
endmodule