module f5_test_7(input in, output reg out);
always @(in)
    out = in;
endmodule