module INV_5 (
	input A,
	output Y
);
	assign Y = !A;
endmodule