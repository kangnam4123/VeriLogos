module U2 (OUT);
   parameter VALUE = 96;
   output [9:0] OUT;
   assign	OUT = VALUE;
endmodule