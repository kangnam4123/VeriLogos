module index___uint16_uint16__uint8_7_3___1(input CLK, input process_CE, input [199:0] inp, output [167:0] process_output);
parameter INSTANCE_NAME="INST";
  assign process_output = (inp[199:32]);
endmodule