module f32_test(output out, input in);
assign out = +in;
endmodule