module sub_7;
   wire pub ;   
   localparam THREE = 3;
endmodule