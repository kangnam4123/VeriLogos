module OR_1
( 
  A, 
  B,
  Z
);
  input A, B;
  output Z;
  assign Z = A|B;
endmodule