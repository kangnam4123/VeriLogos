module GSR_2(output wire GSR);
	assign GSR = 1;
endmodule