module v959751_v465065 #(
 parameter VALUE = 0
) (
 output [31:0] k
);
 assign k = VALUE;
endmodule