module sysgen_constant_118900d9b9 (
  output [(2 - 1):0] op,
  input clk,
  input ce,
  input clr);
  assign op = 2'b11;
endmodule