module JCBUFB1(A, O);
input   A;
output  O;
buf g0(O, A);
endmodule