module GeneratorUnsigned1(out);
	output wire out;
	assign out = 1;
endmodule