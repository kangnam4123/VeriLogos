module sub_40;
   wire pub ;   
endmodule