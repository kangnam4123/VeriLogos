module f1_TECH_AND4(input [3:0] in, output out);
assign out = &in;
endmodule