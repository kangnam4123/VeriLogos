module v2(a, c);
    input [193:0] a;
    output [193:0] c;
    assign c[1:0] = a[187:186];
    assign c[3:2] = 0;
    assign c[5:4] = 0;
    assign c[7:6] = a[189:188];
    assign c[9:8] = 0;
    assign c[11:10] = 0;
    assign c[13:12] = a[191:190];
    assign c[15:14] = 0;
    assign c[17:16] = 0;
    assign c[19:18] = a[185:184];
    assign c[21:20] = 0;
    assign c[23:22] = 0;
    assign c[25:24] = 0;
    assign c[27:26] = a[123:122];
    assign c[29:28] = 0;
    assign c[31:30] = 0;
    assign c[33:32] = a[141:140];
    assign c[35:34] = 0;
    assign c[37:36] = 0;
    assign c[39:38] = a[143:142];
    assign c[41:40] = 0;
    assign c[43:42] = 0;
    assign c[45:44] = a[137:136];
    assign c[47:46] = 0;
    assign c[49:48] = 0;
    assign c[51:50] = a[131:130];
    assign c[53:52] = 0;
    assign c[55:54] = 0;
    assign c[57:56] = a[141:140];
    assign c[59:58] = 0;
    assign c[61:60] = 0;
    assign c[63:62] = a[143:142];
    assign c[65:64] = 0;
    assign c[67:66] = 0;
    assign c[69:68] = a[153:152];
    assign c[71:70] = 0;
    assign c[73:72] = 0;
    assign c[75:74] = a[139:138];
    assign c[77:76] = 0;
    assign c[79:78] = 0;
    assign c[81:80] = a[157:156];
    assign c[83:82] = 0;
    assign c[85:84] = 0;
    assign c[87:86] = a[159:158];
    assign c[89:88] = 0;
    assign c[91:90] = 0;
    assign c[93:92] = a[153:152];
    assign c[95:94] = 0;
    assign c[97:96] = 0;
    assign c[99:98] = a[147:146];
    assign c[101:100] = 0;
    assign c[103:102] = 0;
    assign c[105:104] = a[157:156];
    assign c[107:106] = 0;
    assign c[109:108] = 0;
    assign c[111:110] = a[159:158];
    assign c[113:112] = 0;
    assign c[115:114] = 0;
    assign c[117:116] = a[169:168];
    assign c[119:118] = 0;
    assign c[121:120] = 0;
    assign c[123:122] = a[155:154];
    assign c[125:124] = 0;
    assign c[127:126] = 0;
    assign c[129:128] = a[173:172];
    assign c[131:130] = 0;
    assign c[133:132] = 0;
    assign c[135:134] = a[175:174];
    assign c[137:136] = 0;
    assign c[139:138] = 0;
    assign c[141:140] = a[169:168];
    assign c[143:142] = 0;
    assign c[145:144] = 0;
    assign c[147:146] = a[163:162];
    assign c[149:148] = 0;
    assign c[151:150] = 0;
    assign c[153:152] = a[173:172];
    assign c[155:154] = 0;
    assign c[157:156] = 0;
    assign c[159:158] = a[175:174];
    assign c[161:160] = 0;
    assign c[163:162] = 0;
    assign c[165:164] = a[185:184];
    assign c[167:166] = 0;
    assign c[169:168] = 0;
    assign c[171:170] = a[171:170];
    assign c[173:172] = 0;
    assign c[175:174] = 0;
    assign c[177:176] = a[189:188];
    assign c[179:178] = 0;
    assign c[181:180] = 0;
    assign c[183:182] = a[191:190];
    assign c[185:184] = 0;
    assign c[187:186] = 0;
    assign c[189:188] = a[185:184];
    assign c[191:190] = 0;
    assign c[193:192] = 0;
endmodule