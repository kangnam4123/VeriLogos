module m2014_q4i(
	output out);
 	
	assign out = 1'b0;
	
endmodule