module inverter_nick_yay_2 (input A,
						  output Z);
	assign z = ~A;
endmodule