module MuxN_3(
  input   io_ins_0,
  output  io_out
);
  assign io_out = io_ins_0;
endmodule