module GP_VSS(output OUT);
       assign OUT = 0;
endmodule