module N1Z000( O );     
    output  O;
assign O = 1'b0;
endmodule