module bw_clk_cl_ctu_2xcmp(bw_pll_2x_clk_local ,bw_pll_2xclk );
output		bw_pll_2x_clk_local ;
input		bw_pll_2xclk ;
assign  bw_pll_2x_clk_local =  bw_pll_2xclk;
endmodule