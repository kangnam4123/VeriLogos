module GeneratorSigned1(out);
	output wire signed out;
	assign out = 1;
endmodule