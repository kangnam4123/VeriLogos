module _NOT_(A, Y);
input A;
output Y;
assign Y = ~A;
endmodule