module cyclonev_io_obuf
  (output o, input i, input oe);
   assign o  = i;
   assign oe = oe;
endmodule