module NBUFFX16_1 (INP,Z);
	input INP;
	output Z;
assign Z = INP;
endmodule