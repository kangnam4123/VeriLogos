module v2b9b8c_v9a2a06 (
 input i2,
 input i1,
 input i0,
 output [2:0] o
);
 assign o = {i2, i1, i0};
endmodule