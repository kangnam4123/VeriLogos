module NBUFFX32 (INP,Z);
	input INP;
	output Z;
assign Z = INP;
endmodule