module foobar (clk,d_in, d_out);
input clk;
input  d_in;
output  d_out;
assign d_out = a;
wire  a;
wire  b;
assign a = (b & d_in);
endmodule