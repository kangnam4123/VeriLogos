module bw_clk_cl_ctu_2xcmp_b(bw_pll_2x_clk_local_b ,bw_pll_2xclk_b );
output		bw_pll_2x_clk_local_b ;
input		bw_pll_2xclk_b ;
assign bw_pll_2x_clk_local_b =  bw_pll_2xclk_b;
endmodule