module cp_u4(output wire logic unsigned [7:0] dst,
             input  wire logic unsigned [7:0] src);
  assign dst = src;
endmodule