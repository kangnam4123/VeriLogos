module cycloneiv_io_obuf_1
  (output o, input i, input oe);
   assign o  = i;
   assign oe = oe;
endmodule