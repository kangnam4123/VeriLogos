module BundleBridgeNexus_4(
  input   auto_in,
  output  auto_out_0
);
  assign auto_out_0 = auto_in; 
endmodule