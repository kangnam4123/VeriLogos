module cp_u4s(output wire logic unsigned [3:0] dst,
              input  wire logic unsigned [3:0] src);
  assign dst = src;
endmodule