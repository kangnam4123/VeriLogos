module adder_22 (q,a,b );
input a,b;
output [1:0] q;
assign q =  a  + b;
endmodule