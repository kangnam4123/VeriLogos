module AND2X1_1(A, B, Y);
input A, B;
output Y;
and(Y, A, B);
endmodule