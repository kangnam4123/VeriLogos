module test_27(out);
  output out;
  reg out = 1'b0;
endmodule