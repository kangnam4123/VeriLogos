module Streaminner(
  input   io_input_ctr_done,
  output  io_output_done
);
  assign io_output_done = io_input_ctr_done;
endmodule