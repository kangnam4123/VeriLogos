module packTupleArrays_table__0x0521c798(input CLK, input process_CE, input [335:0] process_input, output [335:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [167:0] unnamedcast2247USEDMULTIPLEcast;assign unnamedcast2247USEDMULTIPLEcast = (process_input[167:0]); 
  wire [167:0] unnamedcast2251USEDMULTIPLEcast;assign unnamedcast2251USEDMULTIPLEcast = (process_input[335:168]); 
  assign process_output = {{({unnamedcast2251USEDMULTIPLEcast[167:160]}),({unnamedcast2247USEDMULTIPLEcast[167:160]})},{({unnamedcast2251USEDMULTIPLEcast[159:152]}),({unnamedcast2247USEDMULTIPLEcast[159:152]})},{({unnamedcast2251USEDMULTIPLEcast[151:144]}),({unnamedcast2247USEDMULTIPLEcast[151:144]})},{({unnamedcast2251USEDMULTIPLEcast[143:136]}),({unnamedcast2247USEDMULTIPLEcast[143:136]})},{({unnamedcast2251USEDMULTIPLEcast[135:128]}),({unnamedcast2247USEDMULTIPLEcast[135:128]})},{({unnamedcast2251USEDMULTIPLEcast[127:120]}),({unnamedcast2247USEDMULTIPLEcast[127:120]})},{({unnamedcast2251USEDMULTIPLEcast[119:112]}),({unnamedcast2247USEDMULTIPLEcast[119:112]})},{({unnamedcast2251USEDMULTIPLEcast[111:104]}),({unnamedcast2247USEDMULTIPLEcast[111:104]})},{({unnamedcast2251USEDMULTIPLEcast[103:96]}),({unnamedcast2247USEDMULTIPLEcast[103:96]})},{({unnamedcast2251USEDMULTIPLEcast[95:88]}),({unnamedcast2247USEDMULTIPLEcast[95:88]})},{({unnamedcast2251USEDMULTIPLEcast[87:80]}),({unnamedcast2247USEDMULTIPLEcast[87:80]})},{({unnamedcast2251USEDMULTIPLEcast[79:72]}),({unnamedcast2247USEDMULTIPLEcast[79:72]})},{({unnamedcast2251USEDMULTIPLEcast[71:64]}),({unnamedcast2247USEDMULTIPLEcast[71:64]})},{({unnamedcast2251USEDMULTIPLEcast[63:56]}),({unnamedcast2247USEDMULTIPLEcast[63:56]})},{({unnamedcast2251USEDMULTIPLEcast[55:48]}),({unnamedcast2247USEDMULTIPLEcast[55:48]})},{({unnamedcast2251USEDMULTIPLEcast[47:40]}),({unnamedcast2247USEDMULTIPLEcast[47:40]})},{({unnamedcast2251USEDMULTIPLEcast[39:32]}),({unnamedcast2247USEDMULTIPLEcast[39:32]})},{({unnamedcast2251USEDMULTIPLEcast[31:24]}),({unnamedcast2247USEDMULTIPLEcast[31:24]})},{({unnamedcast2251USEDMULTIPLEcast[23:16]}),({unnamedcast2247USEDMULTIPLEcast[23:16]})},{({unnamedcast2251USEDMULTIPLEcast[15:8]}),({unnamedcast2247USEDMULTIPLEcast[15:8]})},{({unnamedcast2251USEDMULTIPLEcast[7:0]}),({unnamedcast2247USEDMULTIPLEcast[7:0]})}};
endmodule