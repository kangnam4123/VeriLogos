module vef98b5_v465065 #(
 parameter VALUE = 0
) (
 output [23:0] k
);
 assign k = VALUE-1;
endmodule