module bug27037;
   reg mem[12:2];
   reg [7:0] i;
endmodule