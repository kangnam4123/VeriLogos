module m_3(x);
   output x;
   reg	  \y.z ;
   assign x = \y.z ;
endmodule