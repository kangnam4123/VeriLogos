module fpga_interconnect_1(
    input datain,
    output dataout
);
    assign dataout = datain;
endmodule