module r_USBTYPEC_REV_HIGH(output wire [7:0] reg_0x07);
	assign reg_0x07=8'h00;
endmodule