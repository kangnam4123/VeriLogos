module two (a, b);
   input a, b;
   reg x;
endmodule