module INV_12(output O, input I);
  assign O = !I;
endmodule