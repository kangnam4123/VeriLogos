module f1_test_9(input [1:0] in, output reg [1:0] out);
always @(in)
    out = in;
endmodule