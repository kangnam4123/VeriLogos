module sky130_fd_sc_hvl__lsbuflv2hv_symmetric_2 (
    X,
    A
);
    output X;
    input  A;
    buf buf0 (X     , A              );
endmodule