module FP17_TO_FP16_mgc_in_wire_wait_v1 (ld, vd, d, lz, vz, z);
  parameter integer rscid = 1;
  parameter integer width = 8;
  input ld;
  output vd;
  output [width-1:0] d;
  output lz;
  input vz;
  input [width-1:0] z;
  wire vd;
  wire [width-1:0] d;
  wire lz;
  assign d = z;
  assign lz = ld;
  assign vd = vz;
endmodule