module s1_1(clk, b, so);
input 	clk;
input 	[1:6] b;
output 	[1:4] so;
reg 	[1:4] so;
	always @(posedge clk)
		casex(b)
				6'b000000 :	so=4'he;
				6'b000010 :	so=4'h4;
				6'b000100 :	so=4'hd;
				6'b000110 :	so=4'h1;
				6'b001000 :	so=4'h2;
				6'b001010 :	so=4'hf;
				6'b001100 :	so=4'hb;
				6'b001110 :	so=4'h8;
				6'b010000 :	so=4'h3;
				6'b010010 :	so=4'ha;
				6'b010100 :	so=4'h6;
				6'b010110 :	so=4'hc;
				6'b011000 :	so=4'h5;
				6'b011010 :	so=4'h9;
				6'b011100 :	so=4'h0;
				6'b011110 :	so=4'h7;
				6'b000001 :	so=4'h0;
				6'b000011 :	so=4'hf;
				6'b000101 :	so=4'h7;
				6'b000111 :	so=4'h4;
				6'b001001 :	so=4'he;
				6'b001011 :	so=4'h2;
				6'b001101 :	so=4'hd;
				6'b001111 :	so=4'h1;
				6'b010001 :	so=4'ha;
				6'b010011 :	so=4'h6;
				6'b010101 :	so=4'hc;
				6'b010111 :	so=4'hb;
				6'b011001 :	so=4'h9;
				6'b011011 :	so=4'h5;
				6'b011101 :	so=4'h3;
				6'b011111 :	so=4'h8;
				6'b100000 :	so=4'h4;
				6'b100010 :	so=4'h1;
				6'b100100 :	so=4'he;
				6'b100110 :	so=4'h8;
				6'b101000 :	so=4'hd;
				6'b101010 :	so=4'h6;
				6'b101100 :	so=4'h2;
				6'b101110 :	so=4'hb;
				6'b110000 :	so=4'hf;
				6'b110010 :	so=4'hc;
				6'b110100 :	so=4'h9;
				6'b110110 :	so=4'h7;
				6'b111000 :	so=4'h3;
				6'b111010 :	so=4'ha;
				6'b111100 :	so=4'h5;
				6'b111110 :	so=4'h0;
				6'b100001 :	so=4'hf;
				6'b100011 :	so=4'hc;
				6'b100101 :	so=4'h8;
				6'b100111 :	so=4'h2;
				6'b101001 :	so=4'h4;
				6'b101011 :	so=4'h9;
				6'b101101 :	so=4'h1;
				6'b101111 :	so=4'h7;
				6'b110001 :	so=4'h5;
				6'b110011 :	so=4'hb;
				6'b110101 :	so=4'h3;
				6'b110111 :	so=4'he;
				6'b111001 :	so=4'ha;
				6'b111011 :	so=4'h0;
				6'b111101 :	so=4'h6;
				default         so=4'hd;
			endcase
endmodule