module AND_1(O,A,B);
	input wire A,B;
	output wire O;
	assign O = A*B;
endmodule