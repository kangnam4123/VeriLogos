module cell0(Result0);
output Result0;
assign Result0 = 0;
endmodule