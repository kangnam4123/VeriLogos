module sysgen_constant_07b701207a (
  output [(8 - 1):0] op,
  input clk,
  input ce,
  input clr);
  assign op = 8'b11001000;
endmodule