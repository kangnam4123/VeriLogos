module NBUFFX4_1 (INP,Z);
	input INP;
	output Z;
assign Z = INP;
endmodule