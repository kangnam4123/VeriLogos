module hardcaml_lib_vdd
(
    output o
);
    assign o = 1'b1;
endmodule