module DELLN2X2_1 (INP,Z);
	input INP;
	output Z;
	assign Z  = INP;
endmodule