module OptimizationBarrier_41(
  input  [2:0] io_x,
  output [2:0] io_y
);
  assign io_y = io_x; 
endmodule