module rom (
    dout,
    addr
);
output [7:0] dout;
reg [7:0] dout;
input [6:0] addr;
always @(addr) begin: ROM_READ
    case (addr)
        0: dout = 0;
        1: dout = 8;
        2: dout = 28;
        3: dout = 28;
        4: dout = 28;
        5: dout = 28;
        6: dout = 28;
        7: dout = 8;
        8: dout = 0;
        9: dout = 120;
        10: dout = 14;
        11: dout = 7;
        12: dout = 3;
        13: dout = 1;
        14: dout = 1;
        15: dout = 1;
        16: dout = 0;
        17: dout = 0;
        18: dout = 0;
        19: dout = 24;
        20: dout = 62;
        21: dout = 103;
        22: dout = 65;
        23: dout = 0;
        24: dout = 0;
        25: dout = 0;
        26: dout = 12;
        27: dout = 30;
        28: dout = 63;
        29: dout = 107;
        30: dout = 73;
        31: dout = 8;
        32: dout = 0;
        33: dout = 51;
        34: dout = 102;
        35: dout = 108;
        36: dout = 123;
        37: dout = 119;
        38: dout = 101;
        39: dout = 65;
        40: dout = 0;
        41: dout = 0;
        42: dout = 0;
        43: dout = 6;
        44: dout = 63;
        45: dout = 127;
        46: dout = 59;
        47: dout = 41;
        48: dout = 0;
        49: dout = 59;
        50: dout = 30;
        51: dout = 12;
        52: dout = 8;
        53: dout = 24;
        54: dout = 60;
        55: dout = 110;
        56: dout = 0;
        57: dout = 28;
        58: dout = 94;
        59: dout = 56;
        60: dout = 24;
        61: dout = 60;
        62: dout = 102;
        63: dout = 67;
        64: dout = 0;
        65: dout = 99;
        66: dout = 62;
        67: dout = 93;
        68: dout = 127;
        69: dout = 93;
        70: dout = 62;
        71: dout = 99;
        72: dout = 0;
        73: dout = 8;
        74: dout = 68;
        75: dout = 110;
        76: dout = 127;
        77: dout = 110;
        78: dout = 68;
        79: dout = 8;
        80: dout = 0;
        81: dout = 96;
        82: dout = 120;
        83: dout = 62;
        84: dout = 47;
        85: dout = 41;
        86: dout = 97;
        87: dout = 64;
        88: dout = 0;
        89: dout = 12;
        90: dout = 30;
        91: dout = 8;
        92: dout = 60;
        93: dout = 102;
        94: dout = 65;
        95: dout = 0;
        96: dout = 0;
        97: dout = 30;
        98: dout = 3;
        99: dout = 70;
        100: dout = 92;
        101: dout = 80;
        102: dout = 120;
        103: dout = 63;
        104: dout = 0;
        105: dout = 48;
        106: dout = 88;
        107: dout = 64;
        108: dout = 67;
        109: dout = 70;
        110: dout = 108;
        111: dout = 56;
        112: dout = 0;
        113: dout = 127;
        114: dout = 63;
        115: dout = 3;
        116: dout = 3;
        117: dout = 3;
        118: dout = 3;
        119: dout = 3;
        120: dout = 0;
        121: dout = 65;
        122: dout = 99;
        123: dout = 59;
        124: dout = 63;
        125: dout = 47;
        126: dout = 99;
        default: dout = 67;
    endcase
end
endmodule