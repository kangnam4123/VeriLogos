module BUFD (
	input A,
	output Y
);
	assign Y = A;
endmodule