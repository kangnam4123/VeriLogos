module GSR_1 (input GSRI);
	wire GSRO = GSRI;
endmodule