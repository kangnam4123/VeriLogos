module xlnx_glbl
(
  GSR,
  GTS
);
  output GSR;
  output GTS;
  assign GSR = 0;
  assign GTS = 0;
endmodule