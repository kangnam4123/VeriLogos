module fpu_bufrpt_grp4 (
	in,
	out
);
	input [3:0] in;
	output [3:0] out;
	assign out[3:0] = in[3:0];
endmodule