module empty();
   reg x;
endmodule