module r_VENDOR_ID_HIGH(output wire [7:0] reg_0x01);
	assign reg_0x01=8'h00;
endmodule