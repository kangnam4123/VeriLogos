module logic_0_1 (
    output a
);
  assign a = 0;
endmodule