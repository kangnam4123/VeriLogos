module region_mouse_white(input[10:0] x, input[10:0] y, input[10:0] mx, input[10:0] my, output[3:0] yes);
assign yes = (((y==(my+1))&&((x==(mx+1))||0))||((y==(my+2))&&((x==(mx+1))||(x==(mx+2))||0))||((y==(my+3))&&((x==(mx+1))||(x==(mx+2))||(x==(mx+3))||0))||((y==(my+4))&&((x==(mx+1))||(x==(mx+2))||(x==(mx+3))||(x==(mx+4))||0))||((y==(my+5))&&((x==(mx+1))||(x==(mx+2))||(x==(mx+3))||(x==(mx+4))||(x==(mx+5))||0))||((y==(my+6))&&((x==(mx+1))||(x==(mx+2))||(x==(mx+3))||(x==(mx+4))||(x==(mx+5))||(x==(mx+6))||0))||((y==(my+7))&&((x==(mx+1))||(x==(mx+2))||(x==(mx+3))||(x==(mx+4))||(x==(mx+5))||(x==(mx+6))||(x==(mx+7))||0))||((y==(my+8))&&((x==(mx+1))||(x==(mx+2))||(x==(mx+3))||(x==(mx+4))||(x==(mx+5))||0))||((y==(my+9))&&((x==(mx+1))||(x==(mx+2))||(x==(mx+3))||(x==(mx+4))||(x==(mx+5))||0))||((y==(my+10))&&((x==(mx+1))||(x==(mx+4))||(x==(mx+5))||0))||((y==(my+11))&&((x==(mx+5))||(x==(mx+6))||0))||((y==(my+12))&&((x==(mx+5))||(x==(mx+6))||0))||((y==(my+13))&&((x==(mx+6))||(x==(mx+7))||0))||((y==(my+14))&&((x==(mx+6))||(x==(mx+7))||0))||0) ? 4'b1111 : 4'b0;
endmodule