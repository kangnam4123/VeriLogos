module GP_OBUF(input IN, output OUT);
	assign OUT = IN;
endmodule