module decalper_eb_ot_sdeen_pot_pi_dehcac_xnilix_97
   (In0,
    In1,
    dout);
  input [0:0]In0;
  input [0:0]In1;
  output [1:0]dout;
  wire [0:0]In0;
  wire [0:0]In1;
  assign dout[1] = In1;
  assign dout[0] = In0;
endmodule