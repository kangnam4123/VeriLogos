module xc9500(
  inout wire p34,  
  inout wire p35,
  inout wire p36,  
  inout wire p37,
  inout wire p38,
  inout wire p39,
  inout wire p40,
  inout wire p41,
  inout wire p42,
  inout wire p43,  
  inout wire p44,  
  inout wire p1,   
  inout wire p2,
  inout wire p3,
  inout wire p5,
  inout wire p6,
  inout wire p7,
  inout wire p8,
  inout wire p12,
  inout wire p13,
  inout wire p14,
  inout wire p16,
  inout wire p18,
  inout wire p19,
  inout wire p20,
  inout wire p21,
  inout wire p22,
  inout wire p23,
  inout wire p27,
  inout wire p28,
  inout wire p29,
  inout wire p30,
  inout wire p31,
  inout wire p32,
  inout wire p33  
);
assign p33 = 1'b1;
endmodule