module ANOR6D(A1, A2, A3, A4, A5, A6, O);
input   A1;
input   A2;
input   A3;
input   A4;
input   A5;
input   A6;
output  O;
nor g0(O, A1, A2, A3, A4, A5, A6);
endmodule