module abc9_test008_sub(input a, output b);
assign b = ~a;
endmodule