module INV_13(DATA, RESULT);
input DATA;
output RESULT;
assign RESULT = ~DATA;
endmodule