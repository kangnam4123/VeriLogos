module r_USBPD_REV_VER_HIGH(output wire [7:0] reg_0x09);
	assign reg_0x09=8'h00;
endmodule