module mgc_in_wire (d, z);
  parameter integer rscid = 1;
  parameter integer width = 8;
  output [width-1:0] d;
  input  [width-1:0] z;
  wire   [width-1:0] d;
  assign d = z;
endmodule