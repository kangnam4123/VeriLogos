module s09;
   integer soft; initial soft = 1;
endmodule