module f23_test (out, vout);
output out;
output [7:0] vout;
assign out = 1'b1;
assign vout = 9;
endmodule