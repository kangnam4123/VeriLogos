module N1Z000_1( O );     
    output  O;
assign O = 1'b0;
endmodule