module GP_CLKBUF(input wire IN, output wire OUT);
	assign OUT = IN;
endmodule