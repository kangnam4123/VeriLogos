module inv_1 (input A,
				output Z);
		assign Z = ~A;
	endmodule