module nextReg(X, Y, reset, clk);
   parameter depth=2;
   parameter logDepth=1;
   output Y;
   input X;
   input              clk, reset;
   reg [logDepth:0] count;
   reg                active;
   assign Y = (count == depth) ? 1 : 0;
   always @ (posedge clk) begin
      if (reset == 1) begin
         count <= 0;
         active <= 0;
      end
      else if (X == 1) begin
         active <= 1;
         count <= 1;
      end
      else if (count == depth) begin
         count <= 0;
         active <= 0;
      end
      else if (active)
         count <= count+1;
   end
endmodule