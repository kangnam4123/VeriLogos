module TIELHD (Z);
output Z ;
   buf (Z, 1'B0);
endmodule