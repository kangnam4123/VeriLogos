module cell1(Result0);
output Result0;
assign Result0 = 1;
endmodule