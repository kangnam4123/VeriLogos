module drv1
  (input colSelA,
   output datao
   );
   assign datao = colSelA;
endmodule