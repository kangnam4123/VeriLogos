module glbl_1 ();
    wire GR;
    wire GSR;
    wire GTS;
    wire PRLD;
endmodule