module ham_15_11_encoder (d,c);
	output reg [14:0] c;
	input [10:0] d;
	reg [3:0] p;
	always @(*)
	begin
		p[0]=d[0]^d[1]^d[3]^d[4]^d[6]^d[8]^d[10];
		p[1]=((d[0]^d[2])^(d[3]^d[5]))^((d[6]^d[9])^d[10]);
		p[2]=((d[1]^d[2])^(d[3]^d[7]))^((d[8]^d[9])^d[10]);
		p[3]=((d[4]^d[5])^(d[6]^d[7]))^((d[8]^d[9])^d[10]);
		c[2]=d[0];
		c[4]=d[1];
		c[5]=d[2];
		c[6]=d[3];
		c[8]=d[4];
		c[9]=d[5];
		c[10]=d[6];
		c[11]=d[7];
		c[12]=d[8];
		c[13]=d[9];
		c[14]=d[10];
		c[0]=p[0];
		c[1]=p[1];
		c[3]=p[2];
		c[7]=p[3];
	end
endmodule