module OMUX(L, F, O);
	input wire L;
	input wire F;
	parameter MODE = "";
	output wire O;
	generate
		if ( MODE == "L" )
		begin:SELECT_L
			assign O = L;
		end
		else if ( MODE == "F" )
		begin:SELECT_F
			assign O = F;
		end
		else
		begin
		end
	endgenerate
endmodule