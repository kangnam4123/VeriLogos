module cycloneive_io_obuf_2
  (output o, input i, input oe);
   assign o  = i;
   assign oe = oe;
endmodule