module GND_1(output G);
  assign G = 0;
endmodule