module GP_PWRDET(output reg VDD_LOW);
	initial VDD_LOW = 0;
endmodule