module f7_test_3(output out);
assign out = 1'b0;
endmodule