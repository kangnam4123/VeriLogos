module v3693fc_v465065 #(
 parameter VALUE = 0
) (
 output [4:0] k
);
 assign k = VALUE;
endmodule