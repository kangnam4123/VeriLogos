module submod_1 (b);
   input b;
   reg a;
   initial a = b;
endmodule