module OR2_1 (
	input A, B,
	output Y
);
	assign Y = A | B;
endmodule