module sysgen_constant_1385bcdaec (
  output [(2 - 1):0] op,
  input clk,
  input ce,
  input clr);
  assign op = 2'b11;
endmodule