module WB_SIGN_EXT_8 ( INPUT, OUTPUT );
  input [7:0] INPUT;
  output [31:0] OUTPUT;
  wire   OUTPUT_31;
  assign OUTPUT[31] = OUTPUT_31;
  assign OUTPUT[30] = OUTPUT_31;
  assign OUTPUT[29] = OUTPUT_31;
  assign OUTPUT[28] = OUTPUT_31;
  assign OUTPUT[27] = OUTPUT_31;
  assign OUTPUT[26] = OUTPUT_31;
  assign OUTPUT[25] = OUTPUT_31;
  assign OUTPUT[24] = OUTPUT_31;
  assign OUTPUT[23] = OUTPUT_31;
  assign OUTPUT[22] = OUTPUT_31;
  assign OUTPUT[21] = OUTPUT_31;
  assign OUTPUT[20] = OUTPUT_31;
  assign OUTPUT[19] = OUTPUT_31;
  assign OUTPUT[18] = OUTPUT_31;
  assign OUTPUT[17] = OUTPUT_31;
  assign OUTPUT[16] = OUTPUT_31;
  assign OUTPUT[15] = OUTPUT_31;
  assign OUTPUT[14] = OUTPUT_31;
  assign OUTPUT[13] = OUTPUT_31;
  assign OUTPUT[12] = OUTPUT_31;
  assign OUTPUT[11] = OUTPUT_31;
  assign OUTPUT[10] = OUTPUT_31;
  assign OUTPUT[9] = OUTPUT_31;
  assign OUTPUT[8] = OUTPUT_31;
  assign OUTPUT[7] = OUTPUT_31;
  assign OUTPUT_31 = INPUT[7];
  assign OUTPUT[6] = INPUT[6];
  assign OUTPUT[5] = INPUT[5];
  assign OUTPUT[4] = INPUT[4];
  assign OUTPUT[3] = INPUT[3];
  assign OUTPUT[2] = INPUT[2];
  assign OUTPUT[1] = INPUT[1];
  assign OUTPUT[0] = INPUT[0];
endmodule