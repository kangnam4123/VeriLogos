module LedPattern(
    output wire [('b1000) - ('b1):0] leds);
  assign leds = 'b10010100;
endmodule