module incif_wrapuint32_646_inc2(input CLK, input CE, input [32:0] process_input, output [31:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [31:0] unnamedcast61USEDMULTIPLEcast;assign unnamedcast61USEDMULTIPLEcast = (process_input[31:0]); 
  assign process_output = (((process_input[32]))?((({(unnamedcast61USEDMULTIPLEcast==(32'd646))})?((32'd0)):({(unnamedcast61USEDMULTIPLEcast+(32'd2))}))):(unnamedcast61USEDMULTIPLEcast));
endmodule