module three (a, b, c);
   input a, b, c;
   reg x;
endmodule