module f8_test_1(input in, output out);
assign out = ~in;
endmodule