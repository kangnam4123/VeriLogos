module hdmi_design(clk100, sw, hdmi_rx_scl, hdmi_rx_clk_n, hdmi_rx_clk_p, hdmi_rx_n, hdmi_rx_p, hdmi_tx_hpd, led, debug_pmod, hdmi_rx_cec, hdmi_rx_hpa, hdmi_rx_sda, hdmi_rx_txen, hdmi_tx_cec, hdmi_tx_clk_n, hdmi_tx_clk_p, hdmi_tx_rscl, hdmi_tx_rsda, hdmi_tx_p, hdmi_tx_n, rs232_tx);
  input clk100;
  output [7:0] debug_pmod;
  inout hdmi_rx_cec;
  input hdmi_rx_clk_n;
  input hdmi_rx_clk_p;
  output hdmi_rx_hpa;
  input [2:0] hdmi_rx_n;
  input [2:0] hdmi_rx_p;
  input hdmi_rx_scl;
  inout hdmi_rx_sda;
  output hdmi_rx_txen;
  inout hdmi_tx_cec;
  output hdmi_tx_clk_n;
  output hdmi_tx_clk_p;
  input hdmi_tx_hpd;
  output [2:0] hdmi_tx_n;
  output [2:0] hdmi_tx_p;
  inout hdmi_tx_rscl;
  inout hdmi_tx_rsda;
  output [7:0] led;
  output rs232_tx;
  input [7:0] sw;
  assign hdmi_rx_cec = 1'hz;
  assign hdmi_rx_sda = 1'hz;
  assign hdmi_tx_cec = 1'hz;
  assign hdmi_tx_rscl = 1'hz;
  assign hdmi_tx_rsda = 1'hz;
  assign led = 8'hzz;
  assign debug_pmod = 8'hzz;
  assign hdmi_rx_hpa = 1'hz;
  assign hdmi_rx_txen = 1'hz;
  assign hdmi_tx_clk_n = 1'hz;
  assign hdmi_tx_clk_p = 1'hz;
  assign hdmi_tx_p = 3'hz;
  assign hdmi_tx_n = 3'hz;
  assign rs232_tx = 1'hz;
endmodule