module fpu_bufrpt_grp64 (
	in,
	out
);
	input [63:0] in;
	output [63:0] out;
	assign out[63:0] = in[63:0];
endmodule