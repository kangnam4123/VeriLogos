module v3e6c24_v68c173 (
 output v
);
 assign v = 1'b1;
endmodule