module plane_HV_precomputation (prev_in,A1,A2,B1,B2,shifter1_len,shifter2_len,mux1_sel,mux2_sel,Is7,HV_out);
	input [14:0] prev_in;
	input [7:0] A1,A2,B1,B2;
	input [1:0] shifter1_len,shifter2_len;
	input mux1_sel,mux2_sel;
	input Is7;
	output [14:0] HV_out;
	wire [7:0] neg_A2;
	wire signed [8:0] A1_minus_A2;
	wire signed [11:0] shifter1_out;
	wire [11:0] mux1_out;
	wire [14:0] adder1_out;
	wire [7:0] neg_B2;
	wire signed [8:0] B1_minus_B2;
	wire signed [11:0] shifter2_out;
	wire [9:0] mux2_out;
	wire [9:0] neg_mux2_out;
	wire [11:0] adder2_out;
	assign neg_A2 = ~A2;
	assign A1_minus_A2 = {1'b0,A1} + {1'b1,neg_A2} + 1;	
	assign shifter1_out = A1_minus_A2 <<< shifter1_len;
	assign mux1_out = (mux1_sel == 1'b0)? {{3{A1_minus_A2[8]}},A1_minus_A2}:shifter1_out;
	assign adder1_out = prev_in + {{3{mux1_out[11]}},mux1_out};
	assign neg_B2 = ~B2;
	assign B1_minus_B2 = {1'b0,B1} + {1'b1,neg_B2} + 1;
	assign shifter2_out = B1_minus_B2 <<< shifter2_len;
	assign mux2_out = (mux2_sel == 1'b0)? {B1_minus_B2[8],B1_minus_B2}:{B1_minus_B2,1'b0};
	assign neg_mux2_out = (Is7 == 1'b1)? (~mux2_out + 1):mux2_out;
	assign adder2_out = shifter2_out + {{2{neg_mux2_out[9]}},neg_mux2_out};
	assign HV_out = adder1_out + {{3{adder2_out[11]}},adder2_out};
endmodule