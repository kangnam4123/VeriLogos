module sub_44 (
            input [32:0]  sub_in,
            output [32:0] sub_out);
   assign sub_out = sub_in;
endmodule