module memory_30;
reg [3:0] memory [0:1];
endmodule