module sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_5 (
    X,
    A
);
    output X;
    input  A;
    buf buf0 (X     , A              );
endmodule