module fulladder (a, b, ci, s, co);
  input a, b, ci;
  output co, s;
  wire d;
  assign d = a ^ b;
  assign s = d ^ ci;
  assign co = (b & ~d) | (d & ci);
endmodule