module abc9_test001(input a, output o);
assign o = a;
endmodule