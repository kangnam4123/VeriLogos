module test_25(p);
   output p;
   wire q = 1;
   assign p = q;
endmodule