module cp_s4s(output wire logic signed [3:0] dst,
              input  wire logic signed [3:0] src);
  assign dst = src;
endmodule