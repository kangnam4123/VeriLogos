module f2_test_4(input in, output out);
assign out = ~in;
endmodule