module packTupleArrays_table__0x05765258(input CLK, input process_CE, input [335:0] process_input, output [335:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [167:0] unnamedcast1910USEDMULTIPLEcast;assign unnamedcast1910USEDMULTIPLEcast = (process_input[167:0]); 
  wire [167:0] unnamedcast1914USEDMULTIPLEcast;assign unnamedcast1914USEDMULTIPLEcast = (process_input[335:168]); 
  assign process_output = {{({unnamedcast1914USEDMULTIPLEcast[167:160]}),({unnamedcast1910USEDMULTIPLEcast[167:160]})},{({unnamedcast1914USEDMULTIPLEcast[159:152]}),({unnamedcast1910USEDMULTIPLEcast[159:152]})},{({unnamedcast1914USEDMULTIPLEcast[151:144]}),({unnamedcast1910USEDMULTIPLEcast[151:144]})},{({unnamedcast1914USEDMULTIPLEcast[143:136]}),({unnamedcast1910USEDMULTIPLEcast[143:136]})},{({unnamedcast1914USEDMULTIPLEcast[135:128]}),({unnamedcast1910USEDMULTIPLEcast[135:128]})},{({unnamedcast1914USEDMULTIPLEcast[127:120]}),({unnamedcast1910USEDMULTIPLEcast[127:120]})},{({unnamedcast1914USEDMULTIPLEcast[119:112]}),({unnamedcast1910USEDMULTIPLEcast[119:112]})},{({unnamedcast1914USEDMULTIPLEcast[111:104]}),({unnamedcast1910USEDMULTIPLEcast[111:104]})},{({unnamedcast1914USEDMULTIPLEcast[103:96]}),({unnamedcast1910USEDMULTIPLEcast[103:96]})},{({unnamedcast1914USEDMULTIPLEcast[95:88]}),({unnamedcast1910USEDMULTIPLEcast[95:88]})},{({unnamedcast1914USEDMULTIPLEcast[87:80]}),({unnamedcast1910USEDMULTIPLEcast[87:80]})},{({unnamedcast1914USEDMULTIPLEcast[79:72]}),({unnamedcast1910USEDMULTIPLEcast[79:72]})},{({unnamedcast1914USEDMULTIPLEcast[71:64]}),({unnamedcast1910USEDMULTIPLEcast[71:64]})},{({unnamedcast1914USEDMULTIPLEcast[63:56]}),({unnamedcast1910USEDMULTIPLEcast[63:56]})},{({unnamedcast1914USEDMULTIPLEcast[55:48]}),({unnamedcast1910USEDMULTIPLEcast[55:48]})},{({unnamedcast1914USEDMULTIPLEcast[47:40]}),({unnamedcast1910USEDMULTIPLEcast[47:40]})},{({unnamedcast1914USEDMULTIPLEcast[39:32]}),({unnamedcast1910USEDMULTIPLEcast[39:32]})},{({unnamedcast1914USEDMULTIPLEcast[31:24]}),({unnamedcast1910USEDMULTIPLEcast[31:24]})},{({unnamedcast1914USEDMULTIPLEcast[23:16]}),({unnamedcast1910USEDMULTIPLEcast[23:16]})},{({unnamedcast1914USEDMULTIPLEcast[15:8]}),({unnamedcast1910USEDMULTIPLEcast[15:8]})},{({unnamedcast1914USEDMULTIPLEcast[7:0]}),({unnamedcast1910USEDMULTIPLEcast[7:0]})}};
endmodule