module sum(input  wire [9:0] a, b,
             output wire [9:0] y);
  assign y = a + b;
endmodule