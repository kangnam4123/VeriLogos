module MJBUFDA(A, O);
input   A;
output  O;
buf g0(O, A);
endmodule