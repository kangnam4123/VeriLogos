module IBUF_5(input I, output O);
    assign O = I;
endmodule