module vffc517_v465065 #(
 parameter VALUE = 0
) (
 output [7:0] k
);
 assign k = VALUE;
endmodule