module sky130_fd_sc_lp__busdrivernovlpsleep_2 (
    Z    ,
    A    ,
    TE_B ,
    SLEEP
);
    output Z    ;
    input  A    ;
    input  TE_B ;
    input  SLEEP;
    wire nor_teb_SLEEP;
endmodule