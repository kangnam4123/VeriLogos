module f5_test_5(input in, output out);
assign out = ~in;
endmodule