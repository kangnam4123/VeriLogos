module RAT_xlslice_0_1_1
   (Din,
    Dout);
  input [9:0]Din;
  output [7:0]Dout;
  wire [9:0]Din;
  assign Dout[7:0] = Din[7:0];
endmodule