module test_5;
   parameter foo = 10;
   reg [foo-1:0] bar;
endmodule