module DELLN3X2 (INP,Z);
	input INP;
	output Z;
	assign Z  = INP;
endmodule