module picorv32_regs (
		      input 	    clk, wen,
		      input [5:0]   waddr,
		      input [5:0]   raddr1,
		      input [5:0]   raddr2,
		      input [31:0]  wdata,
		      output [31:0] rdata1,
		      output [31:0] rdata2
		      );
   reg [31:0] 			    regs [0:30];
   always @(posedge clk)
     if (wen) regs[~waddr[4:0]] <= wdata;
   assign rdata1 = regs[~raddr1[4:0]];
   assign rdata2 = regs[~raddr2[4:0]];
endmodule