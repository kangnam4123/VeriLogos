module INVX1(A, Y);
input A;
output Y;
not(Y, A);
endmodule