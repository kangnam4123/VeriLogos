module BUFG_5(output O, input I);
  assign O = I;
endmodule