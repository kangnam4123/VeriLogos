module bsg_counter_clear_up_max_val_p1_init_val_p0
(
  clk_i,
  reset_i,
  clear_i,
  up_i,
  count_o
);
  output [0:0] count_o;
  input clk_i;
  input reset_i;
  input clear_i;
  input up_i;
  wire [0:0] count_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8;
  reg count_o_0_sv2v_reg;
  assign count_o[0] = count_o_0_sv2v_reg;
  always @(posedge clk_i) begin
    if(1'b1) begin
      count_o_0_sv2v_reg <= N8;
    end 
  end
  assign N6 = count_o[0] ^ up_i;
  assign N7 = (N0)? up_i : 
              (N1)? N6 : 1'b0;
  assign N0 = clear_i;
  assign N1 = N5;
  assign N8 = (N2)? 1'b0 : 
              (N3)? N7 : 1'b0;
  assign N2 = reset_i;
  assign N3 = N4;
  assign N4 = ~reset_i;
  assign N5 = ~clear_i;
endmodule