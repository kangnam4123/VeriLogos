module vfebcfe_vb2eccd (
 output q
);
 assign q = 1'b1;
endmodule