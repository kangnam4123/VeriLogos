module OPAD_GTP_VPR (
  input I,
  output O
  );
  assign O = I;
endmodule