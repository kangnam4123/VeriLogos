module z (input i, output oz);
   assign oz = i;
endmodule