module PADIN (output padout, input padin);
   assign padout = padin;
endmodule