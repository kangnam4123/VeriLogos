module r_PD_INTERFACE_REV_HIGH(output wire [7:0] reg_0x0B);
	assign reg_0x0B=8'h00;
endmodule