module GND_2 (output G);
   assign G = 1'b0;
endmodule