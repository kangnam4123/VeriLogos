module constant_9cf45430cd (
  output [(1 - 1):0] op,
  input clk,
  input ce,
  input clr);
  localparam [(1 - 1):0] const_value = 1'b1;
  assign op = 1'b1;
endmodule