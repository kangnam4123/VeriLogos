module fsm_hdlc (
	input clk,
	input reset,
	input in,
	output disc,
	output flag,
	output err);
 	
	parameter [3:0] S0=0, S1=1, S2=2, S3=3, S4=4, S5=5, S6=6, SERR=7, SDISC=8, SFLAG=9;
	reg [3:0] state, next;

	assign disc = state == SDISC;
	assign flag = state == SFLAG;
	assign err = state == SERR;
	
	always @(posedge clk) begin
		case (state)
			S0: state <= in ? S1 : S0;
			S1: state <= in ? S2 : S0;
			S2: state <= in ? S3 : S0;
			S3: state <= in ? S4 : S0;
			S4: state <= in ? S5 : S0;
			S5: state <= in ? S6 : SDISC;
			S6: state <= in ? SERR : SFLAG;
			SERR: state <= in ? SERR : S0;
			SFLAG: state <= in ? S1 : S0;
			SDISC: state <= in ? S1 : S0;
			default: state <= 'x;
		endcase
		
		if (reset) state <= S0;
	end
	
endmodule