module f9_TECH_OR18(input [17:0] in, output out);
assign out = |in;
endmodule