module r_VENDOR_ID_LOW(output wire [7:0] reg_0x00);
	assign reg_0x00=8'h00;
endmodule