module CONNECTNET2(OUT1, OUT2, IN1, IN2);
output OUT1;
output OUT2;
input IN1;
input IN2;
assign OUT1 = IN1;
assign OUT2 = IN2;
endmodule