module v3ba5d0_v465065 #(
 parameter VALUE = 0
) (
 output k
);
 assign k = VALUE;
endmodule