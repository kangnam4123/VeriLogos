module PGAOPV_INVD2PO4 (
  I
 ,ZN
 );
input I ;
output ZN ;
assign ZN = ~I;
endmodule