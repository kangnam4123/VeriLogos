module bw_io_ddr_vref_rptr(in,out,vdd18);
input vdd18;
input [7:0] in;
output [7:0] out;
assign out = in;
endmodule