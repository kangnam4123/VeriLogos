module GP_ABUF(input wire IN, output wire OUT);
	assign OUT = IN;
	parameter BANDWIDTH_KHZ = 1;
endmodule