module U1 (OUT);
   parameter VALUE = -384;
   output [9:0] OUT;
   assign	OUT = VALUE;
endmodule