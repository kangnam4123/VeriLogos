module v3676a0_vd54ca1 (
 input a,
 output q
);
 assign q = ~a;
endmodule