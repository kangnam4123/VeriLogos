module PP1(X, Y, P);
input   X;
input   Y;
output  P;
nor g0(P, X, Y);
endmodule