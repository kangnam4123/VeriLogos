module BundleBridgeNexus_6(
  input   auto_in,
  output  auto_out
);
  assign auto_out = auto_in; 
endmodule