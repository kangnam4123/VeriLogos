module nes_top_X99(a,o);
	input[5:0]  a;
	output reg[7:0]  o;
	always @(a)
	begin
		case(a)
			6'b000000: o = 8'b01101101;
			6'b000001: o = 8'b00100010;
			6'b000010: o = 8'b00000010;
			6'b000011: o = 8'b01000010;
			6'b000100: o = 8'b10000001;
			6'b000101: o = 8'b10100000;
			6'b000110: o = 8'b10100000;
			6'b000111: o = 8'b01100000;
			6'b001000: o = 8'b01000100;
			6'b001001: o = 8'b00001000;
			6'b001010: o = 8'b00001000;
			6'b001011: o = 8'b00000100;
			6'b001100: o = 8'b00000101;
			6'b001101: o = 8'b00000000;
			6'b001110: o = 8'b00000000;
			6'b001111: o = 8'b00000000;
			6'b010000: o = 8'b10110110;
			6'b010001: o = 8'b00001111;
			6'b010010: o = 8'b00100111;
			6'b010011: o = 8'b10000011;
			6'b010100: o = 8'b10100010;
			6'b010101: o = 8'b11100001;
			6'b010110: o = 8'b11000100;
			6'b010111: o = 8'b11001000;
			6'b011000: o = 8'b10001100;
			6'b011001: o = 8'b00010000;
			6'b011010: o = 8'b00010100;
			6'b011011: o = 8'b00010000;
			6'b011100: o = 8'b00010010;
			6'b011101: o = 8'b00000000;
			6'b011110: o = 8'b00000000;
			6'b011111: o = 8'b00000000;
			6'b100000: o = 8'b11111111;
			6'b100001: o = 8'b00110111;
			6'b100010: o = 8'b01010011;
			6'b100011: o = 8'b10110011;
			6'b100100: o = 8'b11101111;
			6'b100101: o = 8'b11101110;
			6'b100110: o = 8'b11101101;
			6'b100111: o = 8'b11110000;
			6'b101000: o = 8'b11110100;
			6'b101001: o = 8'b10011000;
			6'b101010: o = 8'b01011001;
			6'b101011: o = 8'b01011110;
			6'b101100: o = 8'b00011111;
			6'b101101: o = 8'b00000000;
			6'b101110: o = 8'b00000000;
			6'b101111: o = 8'b00000000;
			6'b110000: o = 8'b11111111;
			6'b110001: o = 8'b10111111;
			6'b110010: o = 8'b11011011;
			6'b110011: o = 8'b11011011;
			6'b110100: o = 8'b11111011;
			6'b110101: o = 8'b11111011;
			6'b110110: o = 8'b11110110;
			6'b110111: o = 8'b11111010;
			6'b111000: o = 8'b11111110;
			6'b111001: o = 8'b11111110;
			6'b111010: o = 8'b10111110;
			6'b111011: o = 8'b10111111;
			6'b111100: o = 8'b10011111;
			6'b111101: o = 8'b00000000;
			6'b111110: o = 8'b00000000;
			6'b111111: o = 8'b00000000;
		endcase
	end
endmodule