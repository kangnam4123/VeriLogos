module constant_204e9a8bfd (
  output [(6 - 1):0] op,
  input clk,
  input ce,
  input clr);
  localparam [(6 - 1):0] const_value = 6'b000111;
  assign op = 6'b000111;
endmodule