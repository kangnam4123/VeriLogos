module INVX2(A, Y);
input A;
output Y;
not(Y, A);
endmodule