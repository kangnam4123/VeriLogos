module XOR2X1_1(A, B, Y);
input A, B;
output Y;
xor(Y, A, B);
endmodule