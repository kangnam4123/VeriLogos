module sysgen_constant_61a644b4c8 (
  output [(32 - 1):0] op,
  input clk,
  input ce,
  input clr);
  assign op = 32'b01011111010111100001000000000000;
endmodule