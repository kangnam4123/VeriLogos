module N1Z001_1( O );     
    output  O;
assign O = 1'b1;
endmodule