module f10_TECH_OR5(input [4:0] in, output out);
assign out = |in;
endmodule