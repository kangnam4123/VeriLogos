module BUFX4(A, Y);
input A;
output Y;
buf(Y, A);
endmodule