module f9_TECH_OR4(input [3:0] in, output out);
assign out = |in;
endmodule