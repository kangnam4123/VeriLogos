module RWire0(WHAS, WSET);
   input                    WSET;
   output                   WHAS;
   assign WHAS = WSET;
endmodule