module vio_0_1 (
clk,
probe_out0,
probe_out1,
probe_out2,
probe_out3
);
input clk;
output reg [0 : 0] probe_out0 = 'h0 ;
output reg [0 : 0] probe_out1 = 'h0 ;
output reg [0 : 0] probe_out2 = 'h0 ;
output reg [0 : 0] probe_out3 = 'h0 ;
endmodule