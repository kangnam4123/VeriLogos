module sub_37 (input [3:0] a,
	    output [3:0] z);
   assign z = a;
endmodule