module FP32_MUL_chn_b_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
  assign outsig = in_0;
endmodule