module bsg_buf_width_p1
(
  i,
  o
);
  input [0:0] i;
  output [0:0] o;
  wire [0:0] o;
  assign o[0] = i[0];
endmodule