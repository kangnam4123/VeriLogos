module INVD (
	input A,
	output Y
);
	assign Y = !A;
endmodule