module m2014_q4h(
	input in,
	output out);
 	
	assign out = in;
	
endmodule