module VCC_3(output V);
	assign V = 1;
endmodule