module dec_5to32 (
  input [4:0] a,
  output [31:0] b);  
  and (b[0 ], ~a[4], ~a[3], ~a[2], ~a[1], ~a[0]);
  and (b[1 ], ~a[4], ~a[3], ~a[2], ~a[1],  a[0]);
  and (b[2 ], ~a[4], ~a[3], ~a[2],  a[1], ~a[0]);
  and (b[3 ], ~a[4], ~a[3], ~a[2],  a[1],  a[0]);
  and (b[4 ], ~a[4], ~a[3],  a[2], ~a[1], ~a[0]);
  and (b[5 ], ~a[4], ~a[3],  a[2], ~a[1],  a[0]);
  and (b[6 ], ~a[4], ~a[3],  a[2],  a[1], ~a[0]);
  and (b[7 ], ~a[4], ~a[3],  a[2],  a[1],  a[0]);
  and (b[8 ], ~a[4],  a[3], ~a[2], ~a[1], ~a[0]);
  and (b[9 ], ~a[4],  a[3], ~a[2], ~a[1],  a[0]);
  and (b[10], ~a[4],  a[3], ~a[2],  a[1], ~a[0]);
  and (b[11], ~a[4],  a[3], ~a[2],  a[1],  a[0]);
  and (b[12], ~a[4],  a[3],  a[2], ~a[1], ~a[0]);
  and (b[13], ~a[4],  a[3],  a[2], ~a[1],  a[0]);
  and (b[14], ~a[4],  a[3],  a[2],  a[1], ~a[0]);
  and (b[15], ~a[4],  a[3],  a[2],  a[1],  a[0]);
  and (b[16],  a[4], ~a[3], ~a[2], ~a[1], ~a[0]);
  and (b[17],  a[4], ~a[3], ~a[2], ~a[1],  a[0]);
  and (b[18],  a[4], ~a[3], ~a[2],  a[1], ~a[0]);
  and (b[19],  a[4], ~a[3], ~a[2],  a[1],  a[0]);
  and (b[20],  a[4], ~a[3],  a[2], ~a[1], ~a[0]);
  and (b[21],  a[4], ~a[3],  a[2], ~a[1],  a[0]);
  and (b[22],  a[4], ~a[3],  a[2],  a[1], ~a[0]);
  and (b[23],  a[4], ~a[3],  a[2],  a[1],  a[0]);
  and (b[24],  a[4],  a[3], ~a[2], ~a[1], ~a[0]);
  and (b[25],  a[4],  a[3], ~a[2], ~a[1],  a[0]);
  and (b[26],  a[4],  a[3], ~a[2],  a[1], ~a[0]);
  and (b[27],  a[4],  a[3], ~a[2],  a[1],  a[0]);
  and (b[28],  a[4],  a[3],  a[2], ~a[1], ~a[0]);
  and (b[29],  a[4],  a[3],  a[2], ~a[1],  a[0]);
  and (b[30],  a[4],  a[3],  a[2],  a[1], ~a[0]);
  and (b[31],  a[4],  a[3],  a[2],  a[1],  a[0]);
endmodule