module CARRY_CO_DIRECT_1(input CO, input O, input S, input DI, output OUT);
assign OUT = CO;
endmodule