module hexturnoff (hex6, hex2);
	output [0:6] hex6;
	output [0:6] hex2;
	assign hex6 = 7'b1111111;
	assign hex2 = 7'b1111111;
endmodule