module INC1 #(parameter SIZE = 1) (input in, output [SIZE:0] out);
assign out = in + 1;
endmodule