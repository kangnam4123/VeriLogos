module GP_DAC(input[7:0] DIN, input wire VREF, output reg VOUT);
	initial VOUT = 0;
endmodule