module bsg_mul_csa
     (input x_i
      ,input y_i
      ,input z_i
      ,output c_o
      ,output s_o
      );
     assign {c_o,s_o} = x_i + y_i + z_i;
endmodule