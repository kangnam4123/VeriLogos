module r_PRODUCT_ID_LOW(output wire [7:0] reg_0x02);
	assign reg_0x02=8'h00;
endmodule