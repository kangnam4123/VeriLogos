module GP_INV(input IN, output OUT);
	assign OUT = ~IN;
endmodule