module cp_s4l(output wire logic signed [11:0] dst,
              input  wire logic signed [11:0] src);
  assign dst = src;
endmodule