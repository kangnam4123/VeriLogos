module onewire(input  W_IN, output W_OUT);
  assign W_OUT = W_IN;
endmodule