module r_USBTYPEC_REV_LOW(output wire [7:0] reg_0x06);
	assign reg_0x06=8'h00;
endmodule