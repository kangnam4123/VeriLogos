module glob(fake);
   input fake;
   reg var1;
   reg var2;
endmodule