module logic_0(output a);
    assign a = 0;
endmodule