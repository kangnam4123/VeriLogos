module INVX8(A, Y);
input A;
output Y;
not(Y, A);
endmodule