module VCC(output P);
  assign P = 1;
endmodule