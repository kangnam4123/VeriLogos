module vd4bd04_v9a2a06 (
 input i1,
 input i0,
 output [1:0] o
);
 assign o = {i1, i0};
endmodule