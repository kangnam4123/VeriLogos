module nop(d,q);
input [31:0] d;
output [31:0] q;
  assign q=d;
endmodule