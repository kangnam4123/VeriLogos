module XNOR2X1_1(A, B, Y);
input A, B;
output Y;
xnor(Y, A, B);
endmodule