module hexdisp_eq_2(leds);
	output [0:6] leds;
	assign leds = 7'b1110110; 
endmodule