module _90_lcu_1 (P, G, CI, CO);
	parameter WIDTH = 2;
	input [WIDTH-1:0] P, G;
	input CI;
	output [WIDTH-1:0] CO;
	integer i, j;
	reg [WIDTH-1:0] p, g;
	wire [1023:0] _TECHMAP_DO_ = "proc; opt -fast";
	always @* begin
		p = P;
		g = G;
		g[0] = g[0] | (p[0] & CI);
		for (i = 1; i <= $clog2(WIDTH); i = i+1) begin
			for (j = 2**i - 1; j < WIDTH; j = j + 2**i) begin
				g[j] = g[j] | p[j] & g[j - 2**(i-1)];
				p[j] = p[j] & p[j - 2**(i-1)];
			end
		end
		for (i = $clog2(WIDTH); i > 0; i = i-1) begin
			for (j = 2**i + 2**(i-1) - 1; j < WIDTH; j = j + 2**i) begin
				g[j] = g[j] | p[j] & g[j - 2**(i-1)];
				p[j] = p[j] & p[j - 2**(i-1)];
			end
		end
	end
	assign CO = g;
endmodule