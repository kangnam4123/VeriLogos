module IntXbar(
  input   auto_int_in_0,
  output  auto_int_out_0
);
  assign auto_int_out_0 = auto_int_in_0; 
endmodule