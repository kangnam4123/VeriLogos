module incif_wrapuint32_153615_inc1(input CLK, input CE, input [32:0] process_input, output [31:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [31:0] unnamedcast8525USEDMULTIPLEcast;assign unnamedcast8525USEDMULTIPLEcast = (process_input[31:0]); 
  assign process_output = (((process_input[32]))?((({(unnamedcast8525USEDMULTIPLEcast==(32'd153615))})?((32'd0)):({(unnamedcast8525USEDMULTIPLEcast+(32'd1))}))):(unnamedcast8525USEDMULTIPLEcast));
endmodule