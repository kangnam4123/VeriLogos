module S3(
    input [5:0] B,
    output [3:0] S_B
    );
	 assign S_B =  (B == 0) ? 4'b1010 :
 (B == 1) ? 4'b1101 :
 (B == 2) ? 4'b0 :
 (B == 3) ? 4'b111 :
 (B == 4) ? 4'b1001 :
 (B == 5) ? 4'b0 :
 (B == 6) ? 4'b1110 :
 (B == 7) ? 4'b1001 :
 (B == 8) ? 4'b110 :
 (B == 9) ? 4'b11 :
 (B == 10) ? 4'b11 :
 (B == 11) ? 4'b100 :
 (B == 12) ? 4'b1111 :
 (B == 13) ? 4'b110 :
 (B == 14) ? 4'b101 :
 (B == 15) ? 4'b1010 :
 (B == 16) ? 4'b1 :
 (B == 17) ? 4'b10 :
 (B == 18) ? 4'b1101 :
 (B == 19) ? 4'b1000 :
 (B == 20) ? 4'b1100 :
 (B == 21) ? 4'b101 :
 (B == 22) ? 4'b111 :
 (B == 23) ? 4'b1110 :
 (B == 24) ? 4'b1011 :
 (B == 25) ? 4'b1100 :
 (B == 26) ? 4'b100 :
 (B == 27) ? 4'b1011 :
 (B == 28) ? 4'b10 :
 (B == 29) ? 4'b1111 :
 (B == 30) ? 4'b1000 :
 (B == 31) ? 4'b1 :
 (B == 32) ? 4'b1101 :
 (B == 33) ? 4'b1 :
 (B == 34) ? 4'b110 :
 (B == 35) ? 4'b1010 :
 (B == 36) ? 4'b100 :
 (B == 37) ? 4'b1101 :
 (B == 38) ? 4'b1001 :
 (B == 39) ? 4'b0 :
 (B == 40) ? 4'b1000 :
 (B == 41) ? 4'b110 :
 (B == 42) ? 4'b1111 :
 (B == 43) ? 4'b1001 :
 (B == 44) ? 4'b11 :
 (B == 45) ? 4'b1000 :
 (B == 46) ? 4'b0 :
 (B == 47) ? 4'b111 :
 (B == 48) ? 4'b1011 :
 (B == 49) ? 4'b100 :
 (B == 50) ? 4'b1 :
 (B == 51) ? 4'b1111 :
 (B == 52) ? 4'b10 :
 (B == 53) ? 4'b1110 :
 (B == 54) ? 4'b1100 :
 (B == 55) ? 4'b11 :
 (B == 56) ? 4'b101 :
 (B == 57) ? 4'b1011 :
 (B == 58) ? 4'b1010 :
 (B == 59) ? 4'b101 :
 (B == 60) ? 4'b1110 :
 (B == 61) ? 4'b10 :
 (B == 62) ? 4'b111 : 4'b1100;
endmodule