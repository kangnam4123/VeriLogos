module BUFFER_1 (OUT,IN);
    input IN;
    output OUT;
    buf   ( OUT, IN);
endmodule