module sky130_fd_sc_hdll__nand2b_5 (
    Y  ,
    A_N,
    B
);
    output Y  ;
    input  A_N;
    input  B  ;
    wire not0_out ;
    wire or0_out_Y;
    not not0 (not0_out , B              );
    or  or0  (or0_out_Y, not0_out, A_N  );
    buf buf0 (Y        , or0_out_Y      );
endmodule