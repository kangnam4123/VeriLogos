module ledr(
	input [9:0] buffer,
	output [9:0] lights
	);
	assign lights = buffer;
endmodule