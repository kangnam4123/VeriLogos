module f4_test_5(input [7:0] in, output out);
assign out = ~^in;
endmodule