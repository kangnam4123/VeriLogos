module rom_1 ( input [7:0] addr,output reg [15:0] dout );
always @ (addr)
case (addr)
8'b0000_0000: dout = 16'b0111_0000_0001_0111; 
8'b0000_0001: dout = 16'b1000_0001_0010_0010; 
8'b0000_0010: dout = 16'b1010_0000_0010_0000; 
8'b0000_0011: dout = 16'b1001_0000_0011_0000; 
8'b0000_0100: dout = 16'b0001_0001_0010_0100; 
8'b0000_0101: dout = 16'b0010_0100_0010_0101;  
8'b0000_0110: dout = 16'b1100_0000_0101_0001;  
8'b0000_0111: dout = 16'b1011_0000_0110_0001;  
8'b0000_1000: dout = 16'b0101_0100_0111_0011;  
8'b0000_1001: dout = 16'b0110_0100_1000_0010;  
8'b0000_1010: dout = 16'b0011_0100_0001_1001;  
8'b0000_1011: dout = 16'b0100_0100_0010_1010;  
8'b0000_1100: dout = 16'b1101_0110_0101_0111;  
8'b0000_1101: dout = 16'b0000_0000_0000_0000;  
default:      dout = 16'h0000;
endcase
endmodule