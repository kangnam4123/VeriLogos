module inverter_nick_yay (input A,
						  output Z);
	assign Z = ~A;
endmodule