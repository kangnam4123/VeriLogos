module const_1 (out);
parameter WIDTH=32;
parameter VAL=31;
output [WIDTH-1:0] out;
assign out=VAL;
endmodule