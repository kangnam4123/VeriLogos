module none;
   reg x;
endmodule