module f3_TECH_NAND2(input [1:0] in, output out);
assign out = ~(&in);
endmodule