module Pi(input A, input B, output P);
	assign P = A|B;
endmodule