module f2_TECH_AND5(input [4:0] in, output out);
assign out = &in;
endmodule