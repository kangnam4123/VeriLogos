module sysgen_constant_39c35f37c7 (
  output [(8 - 1):0] op,
  input clk,
  input ce,
  input clr);
  assign op = 8'b11111111;
endmodule